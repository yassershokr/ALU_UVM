package ALU_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "Sequence_item.sv"
    `include "Sequence.sv"
    `include "Sequencer.sv"
    `include "Driver.sv"
    `include "Monitor.sv"
    `include "Coverage_Collector.sv"
    `include "Scoreboard.sv"
    `include "Agent.sv"
    `include "Environment.sv"
    `include "Test.sv"
endpackage: ALU_pkg
